-------------------------------------------------------
--! @file       clkgen.vhd
--! @brief      Clock and reset generator
--! @author     Régis Spadotti (Scalian) 
--! @author     Michel Francis (Scalian)
--! @author     F.Manni (Cnes)
--!
--!-----------------------------------------------------------------------------------------------
--! @copyright  CNES   
--! @verbatim
--! This File is licensed as MIT license
--! Permission is hereby granted, free of charge, to any person obtaining a copy
--! of this software and associated documentation files (the "Software"), to deal
--! in the Software without restriction, including without limitation the rights
--! to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--! copies of the Software, and to permit persons to whom the Software is
--! furnished to do so, subject to the following conditions:
--! 
--! The above copyright notice and this permission notice shall be included in all
--! copies or substantial portions of the Software.
--! 
--! THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--! IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--! FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--! AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--! LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--! OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--! SOFTWARE.
--! @endverbatim
--!
--!-----------------------------------------------------------------------------------------------
--! * Version         : V1.1
--! * Version history : 
--!    * V1 :  2021-03-08 : Scalian : Creation
--!    * V2 :  2021-05-19 : F.Manni (CNES) : 
--!                         * Improve documentation
--! 
--!-----------------------------------------------------------------------------------------------
--! File Creation date : 2021-03-08
--! Project name       : R5 reference Design
--! 
--!-----------------------------------------------------------------------------------------------
--! Softwares             :  
--!     * PC          : Linux Ubuntu 20.04LTS 
--!     * Editor      : Visual studio code 2021-05 + Eclipse 2019-12
--!     * Synthetizer : Nxmap 3.5.0.4 (29th march 2021)
--!     * P&R         : Nxmap 3.5.0.4 (29th march 2021)
--! Automatic VHDL coding :  NO 
--! 
--!-----------------------------------------------------------------------------------------------
--! @details  
--!  
--! @todo provide a detailed description and comments tag for this entity for doxygen
--!
--! Limitations : None
--!
-------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library NX;
use NX.nxPackage.all;

entity clkgen is
port (
   CLK_IN     : in  std_logic; --! external clock on NX140 evalboard : 25 MHz
   RESET      : in  std_logic; --! active high reset 

   CPU_CLK    : out std_logic; --! processor clock : clk vco divided by 4 => 150MHz
   AXI_CLK    : out std_logic; --! processor axi bus frequency : clk vco divided by 20 =>  30MHz
   AXI_CLK_en : out std_logic; --! Axi valid signal for FPGA slaves
                               --! pulse of 1 cpu_clk cycle every axi clk period
                               --! this pulse is centered around axi_clk clock rising edge
                               --! and generated on falling edge of CPU_CLK
   o_CPU_RST_N : out std_logic; --! reset signal active low for cpu domain                           

   APB_CLK    : out std_logic; --! APB clock       :  clk vco divided by 64 : 9.6MH
   o_APB_RST_N : out std_logic; --! reset signal active low for APB domain  

   AHB_CLK    : out std_logic; --! AHB bus clock   : lk vco divided by 80 : 7,5Mhz
   o_AHB_RST_N : out std_logic; --! reset signal active low for AHB domain       

   LOCKED     : out std_logic  --! value 1 when pll is locked
);
end clkgen;

architecture arch of clkgen is
   signal clk_vco         : std_logic; --! vco output signal --600MHZ

   -- first "clock domain" : CPU
   signal clk_vco_div2    : std_logic;    --! clock vco divided by 2 -- 300MHz
   signal clk_vco_div2_div2 : std_logic;  --! clk_vco_div2 divided by 2 by WFG --> 150MHZ
   signal clk_vco_div2_2tap : std_logic;  --! pulse of length of  2 taps of clk_vco_div2 generated by WFG 
   signal clk_vco_div2_div10 : std_logic; --! clk_vco_div2 divided by 10 by WFG --> 30MHZ

   signal rst_pulse_vco_div2 : std_logic; --WFG pulse reset signal (1 period of clk_vco_div2 clock and 1 period before the end of the WFG cycle)
   signal rst_cpu_n : std_logic; --  reset signal 


   -- second clock domain APB
   signal clk_vco_div32   : std_logic;    --! clock vco divided by 32 --  18.75MHZ
   signal clk_vco_div32_div2 : std_logic; --! clock vco divided by 64 => 9.375MHz

   signal rst_pulse_vco_div32 : std_logic; --WFG pulse reset signal (1 period of clk_vco_div32 clock and 1 period before the end of the WFG cycle)
   signal rst_apb_n : std_logic; --  reset signal 

    -- third clock domain : AHB
   signal clk_vco_div8    : std_logic;     --! clock vco divided by 8 --  75Mhz
   signal clk_vco_div8_div_10 : std_logic; --! clock vco divided by 80 --  7,5Mhz

   signal rst_pulse_vco_div8 : std_logic; --WFG pulse reset signal (1 period of clk_vco_div8 clock and 1 period before the end of the WFG cycle)
   signal rst_ahb_n : std_logic; --  reset signal 

   signal sync     : std_logic_vector(4 downto 0); --! synchronization signal for waveform generator patterns
   signal locked_i : std_logic; --! value 1 when PLL is locked

begin

   LOCKED <= locked_i;


 -- # PLL  
   GEN_FREQ : NX_PLL_L
   generic map (
      --! see nxmap libratry guide : chapter 2.4 NX_PLL_L (NG-LARGE) for detailed description
      ref_intdiv => 0,     --! divide input clock by 1 (=> no division) to generate VCO output
      ref_osc_on => '0',   --! use of external clock
      ext_fbk_on => '0',   --! internutilization of internal feedback clock 

      fbk_intdiv   => 10,  --! feedback clock is divided by 10+2 after an intial division by 2
                           --! => clock frequency is then VCO output (or clock input) divided by 24 
      fbk_delay_on => '0', --! no delay for feedback clock
      fbk_delay    => 0,   --! delay set to 0 ()

      clk_outdivp1   => 1, --! clock output p1 divisor : VCO output (=clock input) divided by 2**1 =2           
      clk_outdivp2   => 4, --! clock output p2 divisor : VCO output (=clock input) divided by 2**(4+1) =32       
      clk_outdivo1   => 1, --! clock output o1 divisor : VCO output (=clock input) divided by 2*(1)+3 =5          
      clk_outdivp3o2 => 1  --! clock output p3 and o2 divisor :  VCO output (=clock input) divided by 2*(1)+5 =8           
   )
   port map (
      REF   => CLK_IN,
      FBK   => '0',

      R     => RESET,

      VCO   => clk_vco,
      LDFO  => open,
      REFO  => open,

      DIVO1 => open,
      DIVO2 => clk_vco_div8, 

      DIVP1 => clk_vco_div2,
      DIVP2 => clk_vco_div32, 
      DIVP3 => open,
      OSC   => open,

      PLL_LOCKED => locked_i,
      CAL_LOCKED => open
   );

--------------------------------------------
--
--  # Clock Domain 1 :R5 cluster domain
--  
--
---------------------------------------------

--master WFG (WaveForm Generator) : the one synchronizing output
   busClkEn : NX_WFG_L
   generic map (
      wfg_edge    => '0', -- input clock not inverted
      mode        => '1', -- WFG is used for this clock signal
      pattern_end =>  9,  -- use 10 bits of the patern (if the synchronize signal doesn't reset the pattern before)
      pattern     => "0000011000000000", -- pattern for clock (from left to right bits)
                                         -- this pattern generate a pulse of two clk_vco_div2 tap 
                                         -- at the beginning of the WFG cycle 
      delay_on    => '0'   --no delay
   )
   port map (
      R   => '0',
      SI  => sync(2),
      ZI  => clk_vco_div2,
      RDY => locked_i,
      SO  => sync(2),
      ZO  => clk_vco_div2_2tap);

      AXI_CLK_EN<= clk_vco_div2_2tap;


--"slave1" WFG  synchronized from master 
   WFG_DP1 : NX_WFG_L
     generic map (
       wfg_edge    => '0',-- input clock not inverted
       mode        => '1',-- WFG is used for this clock signal
       pattern_end =>  9, -- use 10 bits of the patern (if the synchronize signal doesn't reset the pattern before)
       pattern     => "1010101010000000", -- pattern for clock (from left to right bits)
                                          -- this pattern create a clock divided by 2
       delay_on    => '0'--no delay
       )
     port map (
       R   => '0',
       SI  => sync(2),
       ZI  => clk_vco_div2,
       RDY => locked_i,
       SO  => sync(0),
       ZO  => clk_vco_div2_div2
       );

       CPU_CLK<=clk_vco_div2_div2;

--"slave2" WFG  synchronized from master
   busClk : NX_WFG_L
     generic map (
       wfg_edge    => '0',-- input clock not inverted
       mode        => '1',-- WFG is used for this clock signal
       pattern_end =>  9, -- use 10 bits of the patern (if the synchronize signal doesn't reset the pattern before)
       pattern     => "0000001111100000",-- pattern for clock (from left to right bits)
                                         -- this pattern divide by 5 the input clock 
       delay_on    => '0'--no delay
       )
     port map (
       R => '0',
       SI => sync(2),
       ZI => clk_vco_div2,
       RDY => locked_i,
       SO => sync(1),
       ZO => clk_vco_div2_div10);

       AXI_CLK<=clk_vco_div2_div10;

--"reset generator  from WFG for CPU domain
-- it uses the fastest clock in the domain
I_CPU_RST : NX_WFG_L
generic map (
  wfg_edge    => '0',-- input clock not inverted
  mode        => '1',-- WFG is used for this clock signal
  pattern_end =>  9, -- use 10 bits of the patern (if the synchronize signal doesn't reset the pattern before)
  pattern     => "0000000110000000",-- pattern for clock (from left to right bits)
                                    -- it provide a pulse of clk_vco_div2 period one clk_vco_div2 period before the end of the WFG cycle 
  delay_on    => '0'--no delay
  )
port map (
  R => '0',
  SI => sync(2),
  ZI => clk_vco_div2,
  RDY => locked_i,
  SO => open,
  ZO => rst_pulse_vco_div2);

  --the reset is released after the rising edge of the fastest clock in the domain
  process(clk_vco_div2_div2,locked_i)
  begin
  if locked_i='0' then
      --PLL not locked => stay in reset
      rst_cpu_n<='0';
  elsif rising_edge(clk_vco_div2_div2) then
      if rst_pulse_vco_div2 ='1' then
         --wait for end of 1st WFG cycle to remove reset
         rst_cpu_n<='1';  
      end if;
   end if;
  end process;
  
  o_CPU_RST_N<=rst_cpu_n; 

--------------------------------------------
--
--  # Clock Domain 2 :APB domain
--  
--
---------------------------------------------
--independant WFG => phase not garanted regarding other WFG (sync input is different)
  WFG_DP2 : NX_WFG_L
   generic map (
      wfg_edge    => '0',-- input clock not inverted
      mode        => '1',-- WFG is used for this clock signal
      pattern_end =>  5, -- use 6 bits of the patern (if the synchronize signal doesn't reset the pattern before)
      pattern     => "1010100000000000",-- pattern for clock (from left to right bits)
                                        -- this pattern divides by two the input clock  
      delay_on    => '0'--no delay
   )
   port map (
      R   => '0',
      SI  => sync(3),
      ZI  => clk_vco_div32,
      RDY => locked_i,
      SO  => sync(3),
      ZO  => clk_vco_div32_div2
   );

   APB_CLK<=clk_vco_div32_div2;


--"reset generator  from WFG for APB domain
I_APB_RST : NX_WFG_L
generic map (
  wfg_edge    => '0',-- input clock not inverted
  mode        => '1',-- WFG is used for this clock signal
  pattern_end =>  5, -- use 10 bits of the patern (if the synchronize signal doesn't reset the pattern before)
  pattern     => "0001100000000000",-- pattern for clock (from left to right bits)
                                    -- it provide a pulse of clk_vco_div2 period one clk_vco_div2 period before the end of the WFG cycle 
  delay_on    => '0'--no delay
  )
port map (
  R => '0',
  SI => sync(3),
  ZI => clk_vco_div32,
  RDY => locked_i,
  SO => open,
  ZO => rst_pulse_vco_div32);

  process(clk_vco_div32_div2,locked_i)
  begin
  if locked_i='0' then
      --PLL not locked => stay in reset
      rst_apb_n<='0';
  elsif rising_edge(clk_vco_div32_div2) then
      if rst_pulse_vco_div32 ='1' then
         --wait for end of 1st WFG cycle to remove reset
         rst_apb_n<='1';  
      end if;
   end if;
  end process;
  o_APB_RST_N<=rst_apb_n;

--------------------------------------------
--
--  Clock Domain 3 : AHB domain
--  
--
---------------------------------------------
--independant WFG => phase not garanted regarding other WFG (sync input is different)
   WFG_DO2 : NX_WFG_L
   generic map (
      wfg_edge    => '0',-- input clock not inverted
      mode        => '1',-- WFG is used for this clock signal
      pattern_end =>  9, -- use 10 bits of the patern (if the synchronize signal doesn't reset the pattern before)
      pattern     => "1110000011000000",-- pattern for clock (from left to right bits)
      delay_on    => '0'--no delay
   )
   port map (
      R   => '0',
      SI  => sync(4),
      ZI  => clk_vco_div8,
      RDY => locked_i,
      SO  => sync(4),
      ZO  => clk_vco_div8_div_10
   );

   AHB_CLK<=clk_vco_div8_div_10;
 
--"reset generator  from WFG for AHB domain
   I_AhB_RST : NX_WFG_L
   generic map (
     wfg_edge    => '0',-- input clock not inverted
     mode        => '1',-- WFG is used for this clock signal
     pattern_end =>  9, -- use 10 bits of the patern (if the synchronize signal doesn't reset the pattern before)
     pattern     => "0000000110000000",-- pattern for clock (from left to right bits)
                                       -- it provide a pulse of clk_vco_div2 period one clk_vco_div2 period before the end of the WFG cycle 
     delay_on    => '0'--no delay
     )
   port map (
     R => '0',
     SI => sync(4),
     ZI => clk_vco_div8,
     RDY => locked_i,
     SO => open,
     ZO => rst_pulse_vco_div8);
   
     process(clk_vco_div8_div_10,locked_i)
     begin
     if locked_i='0' then
         --PLL not locked => stay in reset
         rst_ahb_n<='0';
     elsif rising_edge(clk_vco_div8_div_10) then
         if rst_pulse_vco_div8 ='1' then
            --wait for end of 1st WFG cycle to remove reset
            rst_ahb_n<='1';  
         end if;
      end if;
     end process;
     o_AHB_RST_N<=rst_ahb_n;

end arch;
